LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY decoder_termometrico IS PORT (

	X : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));

END decoder_termometrico;
ARCHITECTURE arc_decoder OF decoder_termometrico IS BEGIN

	S <= "0000000000000001" WHEN X = "0000" ELSE
		"0000000000000011" WHEN X = "0001" ELSE
		"0000000000000111" WHEN X = "0010" ELSE
		"0000000000001111" WHEN X = "0011" ELSE
		"0000000000011111" WHEN X = "0100" ELSE
		"0000000000111111" WHEN X = "0101" ELSE
		"0000000001111111" WHEN X = "0110" ELSE
		"0000000011111111" WHEN X = "0111" ELSE
		"0000000111111111" WHEN X = "1000" ELSE
		"0000001111111111" WHEN X = "1001" ELSE
		"0000011111111111" WHEN X = "1010" ELSE
		"0000111111111111" WHEN X = "1011" ELSE
		"0001111111111111" WHEN X = "1100" ELSE
		"0011111111111111" WHEN X = "1101" ELSE
		"0111111111111111" WHEN X = "1110" ELSE
		"1111111111111111";

END arc_decoder;